// soc_system.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                               //                       clk.clk
		output wire        clock_95_clk,                          //                  clock_95.clk
		input  wire        hps_0_f2h_cold_reset_req_reset_n,      //  hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,     // hps_0_f2h_debug_reset_req.reset_n
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents,  //   hps_0_f2h_stm_hw_events.stm_hwevents
		input  wire        hps_0_f2h_warm_reset_req_reset_n,      //  hps_0_f2h_warm_reset_req.reset_n
		output wire        hps_0_h2f_reset_reset_n,               //           hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK, //              hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,   //                          .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,   //                          .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,   //                          .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,   //                          .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,   //                          .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,   //                          .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,    //                          .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL, //                          .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL, //                          .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK, //                          .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,   //                          .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,   //                          .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,   //                          .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,     //                          .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,     //                          .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,     //                          .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,     //                          .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,     //                          .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,     //                          .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,     //                          .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,      //                          .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,      //                          .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,     //                          .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,      //                          .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,      //                          .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,      //                          .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,      //                          .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,      //                          .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,      //                          .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,      //                          .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,      //                          .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,      //                          .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,      //                          .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,     //                          .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,     //                          .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,     //                          .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,     //                          .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,    //                          .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,   //                          .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,   //                          .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,    //                          .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,     //                          .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,     //                          .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,     //                          .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,     //                          .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,     //                          .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,     //                          .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,  //                          .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,  //                          .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,  //                          .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,  //                          .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,  //                          .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,  //                          .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,  //                          .hps_io_gpio_inst_GPIO61
		output wire [14:0] memory_mem_a,                          //                    memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //                          .mem_ba
		output wire        memory_mem_ck,                         //                          .mem_ck
		output wire        memory_mem_ck_n,                       //                          .mem_ck_n
		output wire        memory_mem_cke,                        //                          .mem_cke
		output wire        memory_mem_cs_n,                       //                          .mem_cs_n
		output wire        memory_mem_ras_n,                      //                          .mem_ras_n
		output wire        memory_mem_cas_n,                      //                          .mem_cas_n
		output wire        memory_mem_we_n,                       //                          .mem_we_n
		output wire        memory_mem_reset_n,                    //                          .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                         //                          .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                        //                          .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                      //                          .mem_dqs_n
		output wire        memory_mem_odt,                        //                          .mem_odt
		output wire [3:0]  memory_mem_dm,                         //                          .mem_dm
		input  wire        memory_oct_rzqin,                      //                          .oct_rzqin
		input  wire [31:0] pio_status_export,                     //                pio_status.export
		input  wire        reset_reset_n                          //                     reset.reset_n
	);

	wire          systolic_array_buffered_0_data_out_valid;                    // systolic_array_buffered_0:data_out_valid -> msgdma_write:st_sink_valid
	wire  [255:0] systolic_array_buffered_0_data_out_data;                     // systolic_array_buffered_0:data_out_data -> msgdma_write:st_sink_data
	wire          systolic_array_buffered_0_data_out_ready;                    // msgdma_write:st_sink_ready -> systolic_array_buffered_0:data_out_ready
	wire          sc_fifo_rhs_out_valid;                                       // sc_fifo_rhs:out_valid -> systolic_array_buffered_0:st_cols_valid
	wire  [255:0] sc_fifo_rhs_out_data;                                        // sc_fifo_rhs:out_data -> systolic_array_buffered_0:st_cols_data
	wire          sc_fifo_rhs_out_ready;                                       // systolic_array_buffered_0:st_cols_ready -> sc_fifo_rhs:out_ready
	wire          sc_fifo_lhs_out_valid;                                       // sc_fifo_lhs:out_valid -> systolic_array_buffered_0:st_rows_valid
	wire  [255:0] sc_fifo_lhs_out_data;                                        // sc_fifo_lhs:out_data -> systolic_array_buffered_0:st_rows_data
	wire          sc_fifo_lhs_out_ready;                                       // systolic_array_buffered_0:st_rows_ready -> sc_fifo_lhs:out_ready
	wire          demux_cols_rows_out0_valid;                                  // demux_cols_rows:out0_valid -> sc_fifo_rhs:in_valid
	wire  [255:0] demux_cols_rows_out0_data;                                   // demux_cols_rows:out0_data -> sc_fifo_rhs:in_data
	wire          demux_cols_rows_out0_ready;                                  // sc_fifo_rhs:in_ready -> demux_cols_rows:out0_ready
	wire          demux_cols_rows_out1_valid;                                  // demux_cols_rows:out1_valid -> sc_fifo_lhs:in_valid
	wire  [255:0] demux_cols_rows_out1_data;                                   // demux_cols_rows:out1_data -> sc_fifo_lhs:in_data
	wire          demux_cols_rows_out1_ready;                                  // sc_fifo_lhs:in_ready -> demux_cols_rows:out1_ready
	wire          msgdma_read_st_source_valid;                                 // msgdma_read:st_source_valid -> demux_cols_rows:in_valid
	wire  [255:0] msgdma_read_st_source_data;                                  // msgdma_read:st_source_data -> demux_cols_rows:in_data
	wire          msgdma_read_st_source_ready;                                 // demux_cols_rows:in_ready -> msgdma_read:st_source_ready
	wire          msgdma_read_st_source_channel;                               // msgdma_read:st_source_channel -> demux_cols_rows:in_channel
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                  // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire    [7:0] hps_0_h2f_axi_master_wstrb;                                  // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                 // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                    // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                 // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                  // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                    // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                 // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                 // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                 // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                 // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire   [63:0] hps_0_h2f_axi_master_wdata;                                  // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                   // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                 // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                 // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                 // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                  // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire   [63:0] hps_0_h2f_axi_master_rdata;                                  // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                 // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                 // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                  // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                  // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                  // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                   // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                    // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                 // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                 // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                 // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire   [31:0] mm_interconnect_0_msgdma_read_csr_readdata;                  // msgdma_read:csr_readdata -> mm_interconnect_0:msgdma_read_csr_readdata
	wire    [2:0] mm_interconnect_0_msgdma_read_csr_address;                   // mm_interconnect_0:msgdma_read_csr_address -> msgdma_read:csr_address
	wire          mm_interconnect_0_msgdma_read_csr_read;                      // mm_interconnect_0:msgdma_read_csr_read -> msgdma_read:csr_read
	wire    [3:0] mm_interconnect_0_msgdma_read_csr_byteenable;                // mm_interconnect_0:msgdma_read_csr_byteenable -> msgdma_read:csr_byteenable
	wire          mm_interconnect_0_msgdma_read_csr_write;                     // mm_interconnect_0:msgdma_read_csr_write -> msgdma_read:csr_write
	wire   [31:0] mm_interconnect_0_msgdma_read_csr_writedata;                 // mm_interconnect_0:msgdma_read_csr_writedata -> msgdma_read:csr_writedata
	wire   [31:0] mm_interconnect_0_msgdma_write_csr_readdata;                 // msgdma_write:csr_readdata -> mm_interconnect_0:msgdma_write_csr_readdata
	wire    [2:0] mm_interconnect_0_msgdma_write_csr_address;                  // mm_interconnect_0:msgdma_write_csr_address -> msgdma_write:csr_address
	wire          mm_interconnect_0_msgdma_write_csr_read;                     // mm_interconnect_0:msgdma_write_csr_read -> msgdma_write:csr_read
	wire    [3:0] mm_interconnect_0_msgdma_write_csr_byteenable;               // mm_interconnect_0:msgdma_write_csr_byteenable -> msgdma_write:csr_byteenable
	wire          mm_interconnect_0_msgdma_write_csr_write;                    // mm_interconnect_0:msgdma_write_csr_write -> msgdma_write:csr_write
	wire   [31:0] mm_interconnect_0_msgdma_write_csr_writedata;                // mm_interconnect_0:msgdma_write_csr_writedata -> msgdma_write:csr_writedata
	wire   [31:0] mm_interconnect_0_systolic_array_buffered_0_csr_readdata;    // systolic_array_buffered_0:csr_readdata -> mm_interconnect_0:systolic_array_buffered_0_csr_readdata
	wire    [7:0] mm_interconnect_0_systolic_array_buffered_0_csr_address;     // mm_interconnect_0:systolic_array_buffered_0_csr_address -> systolic_array_buffered_0:csr_address
	wire          mm_interconnect_0_systolic_array_buffered_0_csr_read;        // mm_interconnect_0:systolic_array_buffered_0_csr_read -> systolic_array_buffered_0:csr_read
	wire          mm_interconnect_0_systolic_array_buffered_0_csr_write;       // mm_interconnect_0:systolic_array_buffered_0_csr_write -> systolic_array_buffered_0:csr_write
	wire   [31:0] mm_interconnect_0_systolic_array_buffered_0_csr_writedata;   // mm_interconnect_0:systolic_array_buffered_0_csr_writedata -> systolic_array_buffered_0:csr_writedata
	wire          mm_interconnect_0_msgdma_read_descriptor_slave_waitrequest;  // msgdma_read:descriptor_slave_waitrequest -> mm_interconnect_0:msgdma_read_descriptor_slave_waitrequest
	wire   [31:0] mm_interconnect_0_msgdma_read_descriptor_slave_byteenable;   // mm_interconnect_0:msgdma_read_descriptor_slave_byteenable -> msgdma_read:descriptor_slave_byteenable
	wire          mm_interconnect_0_msgdma_read_descriptor_slave_write;        // mm_interconnect_0:msgdma_read_descriptor_slave_write -> msgdma_read:descriptor_slave_write
	wire  [255:0] mm_interconnect_0_msgdma_read_descriptor_slave_writedata;    // mm_interconnect_0:msgdma_read_descriptor_slave_writedata -> msgdma_read:descriptor_slave_writedata
	wire          mm_interconnect_0_msgdma_write_descriptor_slave_waitrequest; // msgdma_write:descriptor_slave_waitrequest -> mm_interconnect_0:msgdma_write_descriptor_slave_waitrequest
	wire   [31:0] mm_interconnect_0_msgdma_write_descriptor_slave_byteenable;  // mm_interconnect_0:msgdma_write_descriptor_slave_byteenable -> msgdma_write:descriptor_slave_byteenable
	wire          mm_interconnect_0_msgdma_write_descriptor_slave_write;       // mm_interconnect_0:msgdma_write_descriptor_slave_write -> msgdma_write:descriptor_slave_write
	wire  [255:0] mm_interconnect_0_msgdma_write_descriptor_slave_writedata;   // mm_interconnect_0:msgdma_write_descriptor_slave_writedata -> msgdma_write:descriptor_slave_writedata
	wire          mm_interconnect_0_fifo_instr_in_waitrequest;                 // fifo_instr:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_instr_in_waitrequest
	wire    [0:0] mm_interconnect_0_fifo_instr_in_address;                     // mm_interconnect_0:fifo_instr_in_address -> fifo_instr:avalonmm_write_slave_address
	wire          mm_interconnect_0_fifo_instr_in_write;                       // mm_interconnect_0:fifo_instr_in_write -> fifo_instr:avalonmm_write_slave_write
	wire   [31:0] mm_interconnect_0_fifo_instr_in_writedata;                   // mm_interconnect_0:fifo_instr_in_writedata -> fifo_instr:avalonmm_write_slave_writedata
	wire   [31:0] mm_interconnect_0_pio_0_s1_readdata;                         // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire    [1:0] mm_interconnect_0_pio_0_s1_address;                          // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire  [255:0] msgdma_read_mm_read_readdata;                                // mm_interconnect_1:msgdma_read_mm_read_readdata -> msgdma_read:mm_read_readdata
	wire          msgdma_read_mm_read_waitrequest;                             // mm_interconnect_1:msgdma_read_mm_read_waitrequest -> msgdma_read:mm_read_waitrequest
	wire   [31:0] msgdma_read_mm_read_address;                                 // msgdma_read:mm_read_address -> mm_interconnect_1:msgdma_read_mm_read_address
	wire          msgdma_read_mm_read_read;                                    // msgdma_read:mm_read_read -> mm_interconnect_1:msgdma_read_mm_read_read
	wire   [31:0] msgdma_read_mm_read_byteenable;                              // msgdma_read:mm_read_byteenable -> mm_interconnect_1:msgdma_read_mm_read_byteenable
	wire          msgdma_read_mm_read_readdatavalid;                           // mm_interconnect_1:msgdma_read_mm_read_readdatavalid -> msgdma_read:mm_read_readdatavalid
	wire    [7:0] msgdma_read_mm_read_burstcount;                              // msgdma_read:mm_read_burstcount -> mm_interconnect_1:msgdma_read_mm_read_burstcount
	wire  [255:0] mm_interconnect_1_hps_0_f2h_sdram0_data_readdata;            // hps_0:f2h_sdram0_READDATA -> mm_interconnect_1:hps_0_f2h_sdram0_data_readdata
	wire          mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest;         // hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_1:hps_0_f2h_sdram0_data_waitrequest
	wire   [26:0] mm_interconnect_1_hps_0_f2h_sdram0_data_address;             // mm_interconnect_1:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	wire          mm_interconnect_1_hps_0_f2h_sdram0_data_read;                // mm_interconnect_1:hps_0_f2h_sdram0_data_read -> hps_0:f2h_sdram0_READ
	wire          mm_interconnect_1_hps_0_f2h_sdram0_data_readdatavalid;       // hps_0:f2h_sdram0_READDATAVALID -> mm_interconnect_1:hps_0_f2h_sdram0_data_readdatavalid
	wire    [7:0] mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount;          // mm_interconnect_1:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	wire          msgdma_write_mm_write_waitrequest;                           // mm_interconnect_2:msgdma_write_mm_write_waitrequest -> msgdma_write:mm_write_waitrequest
	wire   [31:0] msgdma_write_mm_write_address;                               // msgdma_write:mm_write_address -> mm_interconnect_2:msgdma_write_mm_write_address
	wire   [31:0] msgdma_write_mm_write_byteenable;                            // msgdma_write:mm_write_byteenable -> mm_interconnect_2:msgdma_write_mm_write_byteenable
	wire          msgdma_write_mm_write_write;                                 // msgdma_write:mm_write_write -> mm_interconnect_2:msgdma_write_mm_write_write
	wire  [255:0] msgdma_write_mm_write_writedata;                             // msgdma_write:mm_write_writedata -> mm_interconnect_2:msgdma_write_mm_write_writedata
	wire    [7:0] msgdma_write_mm_write_burstcount;                            // msgdma_write:mm_write_burstcount -> mm_interconnect_2:msgdma_write_mm_write_burstcount
	wire          mm_interconnect_2_hps_0_f2h_sdram1_data_waitrequest;         // hps_0:f2h_sdram1_WAITREQUEST -> mm_interconnect_2:hps_0_f2h_sdram1_data_waitrequest
	wire   [26:0] mm_interconnect_2_hps_0_f2h_sdram1_data_address;             // mm_interconnect_2:hps_0_f2h_sdram1_data_address -> hps_0:f2h_sdram1_ADDRESS
	wire   [31:0] mm_interconnect_2_hps_0_f2h_sdram1_data_byteenable;          // mm_interconnect_2:hps_0_f2h_sdram1_data_byteenable -> hps_0:f2h_sdram1_BYTEENABLE
	wire          mm_interconnect_2_hps_0_f2h_sdram1_data_write;               // mm_interconnect_2:hps_0_f2h_sdram1_data_write -> hps_0:f2h_sdram1_WRITE
	wire  [255:0] mm_interconnect_2_hps_0_f2h_sdram1_data_writedata;           // mm_interconnect_2:hps_0_f2h_sdram1_data_writedata -> hps_0:f2h_sdram1_WRITEDATA
	wire    [7:0] mm_interconnect_2_hps_0_f2h_sdram1_data_burstcount;          // mm_interconnect_2:hps_0_f2h_sdram1_data_burstcount -> hps_0:f2h_sdram1_BURSTCOUNT
	wire          fifo_instr_out_valid;                                        // fifo_instr:avalonst_source_valid -> avalon_st_adapter:in_0_valid
	wire   [31:0] fifo_instr_out_data;                                         // fifo_instr:avalonst_source_data -> avalon_st_adapter:in_0_data
	wire          fifo_instr_out_ready;                                        // avalon_st_adapter:in_0_ready -> fifo_instr:avalonst_source_ready
	wire          avalon_st_adapter_out_0_valid;                               // avalon_st_adapter:out_0_valid -> systolic_array_buffered_0:st_instr_valid
	wire   [31:0] avalon_st_adapter_out_0_data;                                // avalon_st_adapter:out_0_data -> systolic_array_buffered_0:st_instr_data
	wire          avalon_st_adapter_out_0_ready;                               // systolic_array_buffered_0:st_instr_ready -> avalon_st_adapter:out_0_ready
	wire          rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, demux_cols_rows:reset_n, fifo_instr:reset_n, mm_interconnect_0:msgdma_read_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:msgdma_read_reset_n_reset_bridge_in_reset_reset, mm_interconnect_2:msgdma_write_reset_n_reset_bridge_in_reset_reset, msgdma_read:reset_n_reset_n, msgdma_write:reset_n_reset_n, pio_0:reset_n, sc_fifo_lhs:reset, sc_fifo_rhs:reset, systolic_array_buffered_0:reset_sink_reset]
	wire          rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_f2h_sdram1_data_translator_reset_reset_bridge_in_reset_reset]

	soc_system_clk_95 clk_95 (
		.refclk   (clk_clk),        //  refclk.clk
		.rst      (~reset_reset_n), //   reset.reset
		.outclk_0 (clock_95_clk),   // outclk0.clk
		.locked   ()                // (terminated)
	);

	soc_system_demux_cols_rows demux_cols_rows (
		.clk        (clock_95_clk),                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset), // reset.reset_n
		.in_data    (msgdma_read_st_source_data),      //    in.data
		.in_valid   (msgdma_read_st_source_valid),     //      .valid
		.in_ready   (msgdma_read_st_source_ready),     //      .ready
		.in_channel (msgdma_read_st_source_channel),   //      .channel
		.out0_data  (demux_cols_rows_out0_data),       //  out0.data
		.out0_valid (demux_cols_rows_out0_valid),      //      .valid
		.out0_ready (demux_cols_rows_out0_ready),      //      .ready
		.out1_data  (demux_cols_rows_out1_data),       //  out1.data
		.out1_valid (demux_cols_rows_out1_valid),      //      .valid
		.out1_ready (demux_cols_rows_out1_ready)       //      .ready
	);

	soc_system_fifo_instr fifo_instr (
		.wrclock                          (clock_95_clk),                                //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),             // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_instr_in_writedata),   //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_instr_in_write),       //         .write
		.avalonmm_write_slave_address     (mm_interconnect_0_fifo_instr_in_address),     //         .address
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_instr_in_waitrequest), //         .waitrequest
		.avalonst_source_valid            (fifo_instr_out_valid),                        //      out.valid
		.avalonst_source_data             (fifo_instr_out_data),                         //         .data
		.avalonst_source_ready            (fifo_instr_out_ready)                         //         .ready
	);

	soc_system_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (2)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),                      //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n),                     // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),                      //  f2h_warm_reset_req.reset_n
		.f2h_stm_hwevents         (hps_0_f2h_stm_hw_events_stm_hwevents),                  //   f2h_stm_hw_events.stm_hwevents
		.mem_a                    (memory_mem_a),                                          //              memory.mem_a
		.mem_ba                   (memory_mem_ba),                                         //                    .mem_ba
		.mem_ck                   (memory_mem_ck),                                         //                    .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                       //                    .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                        //                    .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                       //                    .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                      //                    .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                      //                    .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                       //                    .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                    //                    .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                         //                    .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                        //                    .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                      //                    .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                        //                    .mem_odt
		.mem_dm                   (memory_mem_dm),                                         //                    .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                      //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),                 //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),                   //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),                   //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),                   //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),                   //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),                   //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),                   //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),                    //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),                 //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),                 //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),                 //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),                   //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),                   //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),                   //                    .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_hps_io_hps_io_qspi_inst_IO0),                     //                    .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_hps_io_hps_io_qspi_inst_IO1),                     //                    .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_hps_io_hps_io_qspi_inst_IO2),                     //                    .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_hps_io_hps_io_qspi_inst_IO3),                     //                    .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_hps_io_hps_io_qspi_inst_SS0),                     //                    .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_hps_io_hps_io_qspi_inst_CLK),                     //                    .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),                     //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),                      //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),                      //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),                     //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),                      //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),                      //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),                      //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),                      //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),                      //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),                      //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),                      //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),                      //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),                      //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),                      //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),                     //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),                     //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),                     //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),                     //                    .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),                    //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),                   //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),                   //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),                    //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),                     //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),                     //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),                     //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),                     //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),                     //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),                     //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),                  //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),                  //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),                  //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_0_hps_io_hps_io_gpio_inst_GPIO48),                  //                    .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),                  //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),                  //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),                  //                    .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                               //           h2f_reset.reset_n
		.f2h_sdram0_clk           (clock_95_clk),                                          //    f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (mm_interconnect_1_hps_0_f2h_sdram0_data_address),       //     f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount),    //                    .burstcount
		.f2h_sdram0_WAITREQUEST   (mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest),   //                    .waitrequest
		.f2h_sdram0_READDATA      (mm_interconnect_1_hps_0_f2h_sdram0_data_readdata),      //                    .readdata
		.f2h_sdram0_READDATAVALID (mm_interconnect_1_hps_0_f2h_sdram0_data_readdatavalid), //                    .readdatavalid
		.f2h_sdram0_READ          (mm_interconnect_1_hps_0_f2h_sdram0_data_read),          //                    .read
		.f2h_sdram1_clk           (clock_95_clk),                                          //    f2h_sdram1_clock.clk
		.f2h_sdram1_ADDRESS       (mm_interconnect_2_hps_0_f2h_sdram1_data_address),       //     f2h_sdram1_data.address
		.f2h_sdram1_BURSTCOUNT    (mm_interconnect_2_hps_0_f2h_sdram1_data_burstcount),    //                    .burstcount
		.f2h_sdram1_WAITREQUEST   (mm_interconnect_2_hps_0_f2h_sdram1_data_waitrequest),   //                    .waitrequest
		.f2h_sdram1_WRITEDATA     (mm_interconnect_2_hps_0_f2h_sdram1_data_writedata),     //                    .writedata
		.f2h_sdram1_BYTEENABLE    (mm_interconnect_2_hps_0_f2h_sdram1_data_byteenable),    //                    .byteenable
		.f2h_sdram1_WRITE         (mm_interconnect_2_hps_0_f2h_sdram1_data_write),         //                    .write
		.h2f_axi_clk              (clock_95_clk),                                          //       h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),                             //      h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),                           //                    .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),                            //                    .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),                           //                    .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),                          //                    .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),                           //                    .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),                          //                    .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),                           //                    .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),                          //                    .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),                          //                    .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),                              //                    .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),                            //                    .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),                            //                    .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),                            //                    .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),                           //                    .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),                           //                    .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),                              //                    .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),                            //                    .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),                           //                    .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),                           //                    .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),                             //                    .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),                           //                    .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),                            //                    .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),                           //                    .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),                          //                    .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),                           //                    .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),                          //                    .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),                           //                    .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),                          //                    .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),                          //                    .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),                              //                    .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),                            //                    .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),                            //                    .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),                            //                    .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),                           //                    .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready)                            //                    .rready
	);

	soc_system_msgdma_read msgdma_read (
		.mm_read_address              (msgdma_read_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (msgdma_read_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (msgdma_read_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (msgdma_read_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (msgdma_read_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (msgdma_read_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_read_burstcount           (msgdma_read_mm_read_burstcount),                             //                 .burstcount
		.clock_clk                    (clock_95_clk),                                               //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                            //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_msgdma_read_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_msgdma_read_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_msgdma_read_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_msgdma_read_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_msgdma_read_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_msgdma_read_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_msgdma_read_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_msgdma_read_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_msgdma_read_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_msgdma_read_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (),                                                           //          csr_irq.irq
		.st_source_data               (msgdma_read_st_source_data),                                 //        st_source.data
		.st_source_valid              (msgdma_read_st_source_valid),                                //                 .valid
		.st_source_ready              (msgdma_read_st_source_ready),                                //                 .ready
		.st_source_channel            (msgdma_read_st_source_channel)                               //                 .channel
	);

	soc_system_msgdma_write msgdma_write (
		.mm_write_address             (msgdma_write_mm_write_address),                               //         mm_write.address
		.mm_write_write               (msgdma_write_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (msgdma_write_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (msgdma_write_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (msgdma_write_mm_write_waitrequest),                           //                 .waitrequest
		.mm_write_burstcount          (msgdma_write_mm_write_burstcount),                            //                 .burstcount
		.clock_clk                    (clock_95_clk),                                                //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                             //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_msgdma_write_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_msgdma_write_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_msgdma_write_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_msgdma_write_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_msgdma_write_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_msgdma_write_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_msgdma_write_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_msgdma_write_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_msgdma_write_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_msgdma_write_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (),                                                            //          csr_irq.irq
		.st_sink_data                 (systolic_array_buffered_0_data_out_data),                     //          st_sink.data
		.st_sink_valid                (systolic_array_buffered_0_data_out_valid),                    //                 .valid
		.st_sink_ready                (systolic_array_buffered_0_data_out_ready)                     //                 .ready
	);

	soc_system_pio_0 pio_0 (
		.clk      (clock_95_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_0_s1_readdata), //                    .readdata
		.in_port  (pio_status_export)                    // external_connection.export
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (32),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (32),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sc_fifo_lhs (
		.clk               (clock_95_clk),                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),       // clk_reset.reset
		.in_data           (demux_cols_rows_out1_data),            //        in.data
		.in_valid          (demux_cols_rows_out1_valid),           //          .valid
		.in_ready          (demux_cols_rows_out1_ready),           //          .ready
		.out_data          (sc_fifo_lhs_out_data),                 //       out.data
		.out_valid         (sc_fifo_lhs_out_valid),                //          .valid
		.out_ready         (sc_fifo_lhs_out_ready),                //          .ready
		.csr_address       (2'b00),                                // (terminated)
		.csr_read          (1'b0),                                 // (terminated)
		.csr_write         (1'b0),                                 // (terminated)
		.csr_readdata      (),                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
		.almost_full_data  (),                                     // (terminated)
		.almost_empty_data (),                                     // (terminated)
		.in_startofpacket  (1'b0),                                 // (terminated)
		.in_endofpacket    (1'b0),                                 // (terminated)
		.out_startofpacket (),                                     // (terminated)
		.out_endofpacket   (),                                     // (terminated)
		.in_empty          (1'b0),                                 // (terminated)
		.out_empty         (),                                     // (terminated)
		.in_error          (1'b0),                                 // (terminated)
		.out_error         (),                                     // (terminated)
		.in_channel        (1'b0),                                 // (terminated)
		.out_channel       ()                                      // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (32),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (32),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sc_fifo_rhs (
		.clk               (clock_95_clk),                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),       // clk_reset.reset
		.in_data           (demux_cols_rows_out0_data),            //        in.data
		.in_valid          (demux_cols_rows_out0_valid),           //          .valid
		.in_ready          (demux_cols_rows_out0_ready),           //          .ready
		.out_data          (sc_fifo_rhs_out_data),                 //       out.data
		.out_valid         (sc_fifo_rhs_out_valid),                //          .valid
		.out_ready         (sc_fifo_rhs_out_ready),                //          .ready
		.csr_address       (2'b00),                                // (terminated)
		.csr_read          (1'b0),                                 // (terminated)
		.csr_write         (1'b0),                                 // (terminated)
		.csr_readdata      (),                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
		.almost_full_data  (),                                     // (terminated)
		.almost_empty_data (),                                     // (terminated)
		.in_startofpacket  (1'b0),                                 // (terminated)
		.in_endofpacket    (1'b0),                                 // (terminated)
		.out_startofpacket (),                                     // (terminated)
		.out_endofpacket   (),                                     // (terminated)
		.in_empty          (1'b0),                                 // (terminated)
		.out_empty         (),                                     // (terminated)
		.in_error          (1'b0),                                 // (terminated)
		.out_error         (),                                     // (terminated)
		.in_channel        (1'b0),                                 // (terminated)
		.out_channel       ()                                      // (terminated)
	);

	systolic_array_top systolic_array_buffered_0 (
		.csr_address      (mm_interconnect_0_systolic_array_buffered_0_csr_address),   //        csr.address
		.csr_write        (mm_interconnect_0_systolic_array_buffered_0_csr_write),     //           .write
		.csr_writedata    (mm_interconnect_0_systolic_array_buffered_0_csr_writedata), //           .writedata
		.csr_readdata     (mm_interconnect_0_systolic_array_buffered_0_csr_readdata),  //           .readdata
		.csr_read         (mm_interconnect_0_systolic_array_buffered_0_csr_read),      //           .read
		.data_out_data    (systolic_array_buffered_0_data_out_data),                   //   data_out.data
		.data_out_ready   (systolic_array_buffered_0_data_out_ready),                  //           .ready
		.data_out_valid   (systolic_array_buffered_0_data_out_valid),                  //           .valid
		.reset_sink_reset (rst_controller_reset_out_reset),                            // reset_sink.reset
		.clock_sink       (clock_95_clk),                                              // clock_sink.clk
		.st_rows_data     (sc_fifo_lhs_out_data),                                      //    st_rows.data
		.st_rows_ready    (sc_fifo_lhs_out_ready),                                     //           .ready
		.st_rows_valid    (sc_fifo_lhs_out_valid),                                     //           .valid
		.st_cols_data     (sc_fifo_rhs_out_data),                                      //    st_cols.data
		.st_cols_ready    (sc_fifo_rhs_out_ready),                                     //           .ready
		.st_cols_valid    (sc_fifo_rhs_out_valid),                                     //           .valid
		.st_instr_ready   (avalon_st_adapter_out_0_ready),                             //   st_instr.ready
		.st_instr_valid   (avalon_st_adapter_out_0_valid),                             //           .valid
		.st_instr_data    (avalon_st_adapter_out_0_data)                               //           .data
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                   //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                                 //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                  //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                                 //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                                //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                                 //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                                //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                                 //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                                //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                                //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                    //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                  //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                  //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                  //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                                 //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                                 //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                    //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                  //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                                 //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                                 //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                   //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                                 //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                  //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                                 //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                                //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                                 //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                                //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                                 //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                                //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                                //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                    //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                  //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                  //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                  //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                                 //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                                 //                                                           .rready
		.clock_bridge_0_out_clk_clk                                       (clock_95_clk),                                                //                                     clock_bridge_0_out_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.msgdma_read_reset_n_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                              //                  msgdma_read_reset_n_reset_bridge_in_reset.reset
		.fifo_instr_in_address                                            (mm_interconnect_0_fifo_instr_in_address),                     //                                              fifo_instr_in.address
		.fifo_instr_in_write                                              (mm_interconnect_0_fifo_instr_in_write),                       //                                                           .write
		.fifo_instr_in_writedata                                          (mm_interconnect_0_fifo_instr_in_writedata),                   //                                                           .writedata
		.fifo_instr_in_waitrequest                                        (mm_interconnect_0_fifo_instr_in_waitrequest),                 //                                                           .waitrequest
		.msgdma_read_csr_address                                          (mm_interconnect_0_msgdma_read_csr_address),                   //                                            msgdma_read_csr.address
		.msgdma_read_csr_write                                            (mm_interconnect_0_msgdma_read_csr_write),                     //                                                           .write
		.msgdma_read_csr_read                                             (mm_interconnect_0_msgdma_read_csr_read),                      //                                                           .read
		.msgdma_read_csr_readdata                                         (mm_interconnect_0_msgdma_read_csr_readdata),                  //                                                           .readdata
		.msgdma_read_csr_writedata                                        (mm_interconnect_0_msgdma_read_csr_writedata),                 //                                                           .writedata
		.msgdma_read_csr_byteenable                                       (mm_interconnect_0_msgdma_read_csr_byteenable),                //                                                           .byteenable
		.msgdma_read_descriptor_slave_write                               (mm_interconnect_0_msgdma_read_descriptor_slave_write),        //                               msgdma_read_descriptor_slave.write
		.msgdma_read_descriptor_slave_writedata                           (mm_interconnect_0_msgdma_read_descriptor_slave_writedata),    //                                                           .writedata
		.msgdma_read_descriptor_slave_byteenable                          (mm_interconnect_0_msgdma_read_descriptor_slave_byteenable),   //                                                           .byteenable
		.msgdma_read_descriptor_slave_waitrequest                         (mm_interconnect_0_msgdma_read_descriptor_slave_waitrequest),  //                                                           .waitrequest
		.msgdma_write_csr_address                                         (mm_interconnect_0_msgdma_write_csr_address),                  //                                           msgdma_write_csr.address
		.msgdma_write_csr_write                                           (mm_interconnect_0_msgdma_write_csr_write),                    //                                                           .write
		.msgdma_write_csr_read                                            (mm_interconnect_0_msgdma_write_csr_read),                     //                                                           .read
		.msgdma_write_csr_readdata                                        (mm_interconnect_0_msgdma_write_csr_readdata),                 //                                                           .readdata
		.msgdma_write_csr_writedata                                       (mm_interconnect_0_msgdma_write_csr_writedata),                //                                                           .writedata
		.msgdma_write_csr_byteenable                                      (mm_interconnect_0_msgdma_write_csr_byteenable),               //                                                           .byteenable
		.msgdma_write_descriptor_slave_write                              (mm_interconnect_0_msgdma_write_descriptor_slave_write),       //                              msgdma_write_descriptor_slave.write
		.msgdma_write_descriptor_slave_writedata                          (mm_interconnect_0_msgdma_write_descriptor_slave_writedata),   //                                                           .writedata
		.msgdma_write_descriptor_slave_byteenable                         (mm_interconnect_0_msgdma_write_descriptor_slave_byteenable),  //                                                           .byteenable
		.msgdma_write_descriptor_slave_waitrequest                        (mm_interconnect_0_msgdma_write_descriptor_slave_waitrequest), //                                                           .waitrequest
		.pio_0_s1_address                                                 (mm_interconnect_0_pio_0_s1_address),                          //                                                   pio_0_s1.address
		.pio_0_s1_readdata                                                (mm_interconnect_0_pio_0_s1_readdata),                         //                                                           .readdata
		.systolic_array_buffered_0_csr_address                            (mm_interconnect_0_systolic_array_buffered_0_csr_address),     //                              systolic_array_buffered_0_csr.address
		.systolic_array_buffered_0_csr_write                              (mm_interconnect_0_systolic_array_buffered_0_csr_write),       //                                                           .write
		.systolic_array_buffered_0_csr_read                               (mm_interconnect_0_systolic_array_buffered_0_csr_read),        //                                                           .read
		.systolic_array_buffered_0_csr_readdata                           (mm_interconnect_0_systolic_array_buffered_0_csr_readdata),    //                                                           .readdata
		.systolic_array_buffered_0_csr_writedata                          (mm_interconnect_0_systolic_array_buffered_0_csr_writedata)    //                                                           .writedata
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.clock_bridge_0_out_clk_clk                                         (clock_95_clk),                                          //                                       clock_bridge_0_out_clk.clk
		.hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.msgdma_read_reset_n_reset_bridge_in_reset_reset                    (rst_controller_reset_out_reset),                        //                    msgdma_read_reset_n_reset_bridge_in_reset.reset
		.msgdma_read_mm_read_address                                        (msgdma_read_mm_read_address),                           //                                          msgdma_read_mm_read.address
		.msgdma_read_mm_read_waitrequest                                    (msgdma_read_mm_read_waitrequest),                       //                                                             .waitrequest
		.msgdma_read_mm_read_burstcount                                     (msgdma_read_mm_read_burstcount),                        //                                                             .burstcount
		.msgdma_read_mm_read_byteenable                                     (msgdma_read_mm_read_byteenable),                        //                                                             .byteenable
		.msgdma_read_mm_read_read                                           (msgdma_read_mm_read_read),                              //                                                             .read
		.msgdma_read_mm_read_readdata                                       (msgdma_read_mm_read_readdata),                          //                                                             .readdata
		.msgdma_read_mm_read_readdatavalid                                  (msgdma_read_mm_read_readdatavalid),                     //                                                             .readdatavalid
		.hps_0_f2h_sdram0_data_address                                      (mm_interconnect_1_hps_0_f2h_sdram0_data_address),       //                                        hps_0_f2h_sdram0_data.address
		.hps_0_f2h_sdram0_data_read                                         (mm_interconnect_1_hps_0_f2h_sdram0_data_read),          //                                                             .read
		.hps_0_f2h_sdram0_data_readdata                                     (mm_interconnect_1_hps_0_f2h_sdram0_data_readdata),      //                                                             .readdata
		.hps_0_f2h_sdram0_data_burstcount                                   (mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount),    //                                                             .burstcount
		.hps_0_f2h_sdram0_data_readdatavalid                                (mm_interconnect_1_hps_0_f2h_sdram0_data_readdatavalid), //                                                             .readdatavalid
		.hps_0_f2h_sdram0_data_waitrequest                                  (mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest)    //                                                             .waitrequest
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.clock_bridge_0_out_clk_clk                                         (clock_95_clk),                                        //                                       clock_bridge_0_out_clk.clk
		.hps_0_f2h_sdram1_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                  // hps_0_f2h_sdram1_data_translator_reset_reset_bridge_in_reset.reset
		.msgdma_write_reset_n_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                      //                   msgdma_write_reset_n_reset_bridge_in_reset.reset
		.msgdma_write_mm_write_address                                      (msgdma_write_mm_write_address),                       //                                        msgdma_write_mm_write.address
		.msgdma_write_mm_write_waitrequest                                  (msgdma_write_mm_write_waitrequest),                   //                                                             .waitrequest
		.msgdma_write_mm_write_burstcount                                   (msgdma_write_mm_write_burstcount),                    //                                                             .burstcount
		.msgdma_write_mm_write_byteenable                                   (msgdma_write_mm_write_byteenable),                    //                                                             .byteenable
		.msgdma_write_mm_write_write                                        (msgdma_write_mm_write_write),                         //                                                             .write
		.msgdma_write_mm_write_writedata                                    (msgdma_write_mm_write_writedata),                     //                                                             .writedata
		.hps_0_f2h_sdram1_data_address                                      (mm_interconnect_2_hps_0_f2h_sdram1_data_address),     //                                        hps_0_f2h_sdram1_data.address
		.hps_0_f2h_sdram1_data_write                                        (mm_interconnect_2_hps_0_f2h_sdram1_data_write),       //                                                             .write
		.hps_0_f2h_sdram1_data_writedata                                    (mm_interconnect_2_hps_0_f2h_sdram1_data_writedata),   //                                                             .writedata
		.hps_0_f2h_sdram1_data_burstcount                                   (mm_interconnect_2_hps_0_f2h_sdram1_data_burstcount),  //                                                             .burstcount
		.hps_0_f2h_sdram1_data_byteenable                                   (mm_interconnect_2_hps_0_f2h_sdram1_data_byteenable),  //                                                             .byteenable
		.hps_0_f2h_sdram1_data_waitrequest                                  (mm_interconnect_2_hps_0_f2h_sdram1_data_waitrequest)  //                                                             .waitrequest
	);

	soc_system_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (0),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk   (clock_95_clk),                   // in_clk_0.clk
		.in_rst_0_reset (rst_controller_reset_out_reset), // in_rst_0.reset
		.in_0_data      (fifo_instr_out_data),            //     in_0.data
		.in_0_valid     (fifo_instr_out_valid),           //         .valid
		.in_0_ready     (fifo_instr_out_ready),           //         .ready
		.out_0_data     (avalon_st_adapter_out_0_data),   //    out_0.data
		.out_0_valid    (avalon_st_adapter_out_0_valid),  //         .valid
		.out_0_ready    (avalon_st_adapter_out_0_ready)   //         .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clock_95_clk),                   //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clock_95_clk),                       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
